module top ()

endmodule